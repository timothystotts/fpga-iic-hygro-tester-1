
localparam [0:0] OP_NONE = 0;
localparam [0:0] OP_POLL_HYGRO = 1;

localparam [2:0] DISP_NONE = 0;
localparam [2:0] DISP_BOTH_CELCIUS = 1;
localparam [2:0] DISP_BOTH_FARH = 2;
localparam [2:0] DISP_ONLY_TEMP_C = 3;
localparam [2:0] DISP_ONLY_TEMP_F = 4;
localparam [2:0] DISP_ONLY_HUMID = 5;
localparam [2:0] DISP_UNKNOWN_A = 6;
localparam [2:0] DISP_UNKNOWN_B = 7;
